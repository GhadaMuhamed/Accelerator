LIBRARY IEEE;
USE IEEE.std_logic_1164.all;

ENTITY mux_8 IS  
Generic (n : integer :=5);
PORT (
IN1,IN2,IN3,IN4,IN5,IN6: IN STD_LOGIC_VECTOR(n-1 DOWNTO 0);
SEl:IN STD_LOGIC_VECTOR(2 DOWNTO 0);
OUT1:OUT  STD_LOGIC_VECTOR(n-1 DOWNTO 0)
);    
END ENTITY mux_8;


ARCHITECTURE ArchMux8 OF mux_8 IS
BEGIN
OUT1 <= IN1 WHEN SEl="000"
ELSE IN2 WHEN SEL="001"
ELSE IN3 WHEN SEL="010"
ELSE IN4 WHEN SEL="011"
ELSE IN5 WHEN SEL="100"
ELSE IN6;
END ArchMux8;
