

LIBRARY IEEE;
USE IEEE.std_logic_1164.all;

ENTITY mux IS  
Generic (n : integer :=17);
PORT (
IN1,IN2,IN3: IN STD_LOGIC_VECTOR(n-1 DOWNTO 0);
SEl:IN STD_LOGIC_VECTOR(1 DOWNTO 0);
OUT1:OUT  STD_LOGIC_VECTOR(n-1 DOWNTO 0)
);    
END ENTITY mux;


ARCHITECTURE ArchMux OF mux IS
BEGIN
OUT1 <= IN1 WHEN SEl="00" OR SEl="01"
ELSE IN2 WHEN SEl="10" 
ELSE IN3 WHEN SEl="11" ;
END ArchMux;