LIBRARY IEEE;
USE IEEE.std_logic_1164.all;

ENTITY pcmux IS  
Generic (n : integer :=17);
PORT (
IN1,IN2,IN3,IN4,IN5,IN6: IN STD_LOGIC_VECTOR(n-1 DOWNTO 0);
SEl:IN STD_LOGIC_VECTOR(2 DOWNTO 0);
OUT1:OUT  STD_LOGIC_VECTOR(n-1 DOWNTO 0)
);    
END ENTITY pcmux;


ARCHITECTURE ArchMux OF pcmux IS
BEGIN
OUT1 <= IN1 WHEN SEl="111" OR SEl="110" 
ELSE IN2 WHEN SEl="101"
ELSE IN3 WHEN SEl="100"
ELSE IN4 WHEN SEl="011"
ELSE IN5 WHEN SEl="010"
ELSE IN6 WHEN SEl="001" OR SEl="000" ;
END ArchMux;